module window

#include <SFML/Window/WindowHandle.h>
