module window

#include <SFML/Window/Types.h>

struct C.sfContext {
}

// Context
pub type Context = C.sfContext

struct C.sfCursor {
}

// Cursor
pub type Cursor = C.sfCursor

struct C.sfWindow {
}

// Window
pub type Window = C.sfWindow
