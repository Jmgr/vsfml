module audio

#include <SFML/Audio/Types.h>

struct C.sfMusic {
}

// Music
pub type Music = C.sfMusic

struct C.sfSound {
}

// Sound
pub type Sound = C.sfSound

struct C.sfSoundBuffer {
}

// SoundBuffer
pub type SoundBuffer = C.sfSoundBuffer

struct C.sfSoundBufferRecorder {
}

// SoundBufferRecorder
pub type SoundBufferRecorder = C.sfSoundBufferRecorder

struct C.sfSoundRecorder {
}

// SoundRecorder
pub type SoundRecorder = C.sfSoundRecorder

struct C.sfSoundStream {
}

// SoundStream
pub type SoundStream = C.sfSoundStream
