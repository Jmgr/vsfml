module window

#include <SFML/Window/Export.h>
