module network

#include <SFML/Network/Types.h>

struct C.sfFtpDirectoryResponse {
}

// FtpDirectoryResponse
pub type FtpDirectoryResponse = C.sfFtpDirectoryResponse

struct C.sfFtpListingResponse {
}

// FtpListingResponse
pub type FtpListingResponse = C.sfFtpListingResponse

struct C.sfFtpResponse {
}

// FtpResponse
pub type FtpResponse = C.sfFtpResponse

struct C.sfFtp {
}

// Ftp
pub type Ftp = C.sfFtp

struct C.sfHttpRequest {
}

// HttpRequest
pub type HttpRequest = C.sfHttpRequest

struct C.sfHttpResponse {
}

// HttpResponse
pub type HttpResponse = C.sfHttpResponse

struct C.sfHttp {
}

// Http
pub type Http = C.sfHttp

struct C.sfPacket {
}

// Packet
pub type Packet = C.sfPacket

struct C.sfSocketSelector {
}

// SocketSelector
pub type SocketSelector = C.sfSocketSelector

struct C.sfTcpListener {
}

// TcpListener
pub type TcpListener = C.sfTcpListener

struct C.sfTcpSocket {
}

// TcpSocket
pub type TcpSocket = C.sfTcpSocket

struct C.sfUdpSocket {
}

// UdpSocket
pub type UdpSocket = C.sfUdpSocket
