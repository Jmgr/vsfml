// system: base module of SFML, defining various utilities
module system

#flag -lcsfml-system
