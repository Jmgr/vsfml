// audio: sounds, streaming (musics or custom sources), recording, spatialization
module audio

#flag -lcsfml-audio
