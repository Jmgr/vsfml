module system

#include <SFML/System/Types.h>

struct C.sfClock {
}

// Clock
pub type Clock = C.sfClock

struct C.sfMutex {
}

// Mutex
pub type Mutex = C.sfMutex

struct C.sfThread {
}

// Thread
pub type Thread = C.sfThread
