// graphics: 2D graphics module: sprites, text, shapes, ...
module graphics

#flag -I @VROOT/graphics/c
#flag @VROOT/graphics/c/graphics.c
#include "graphics.h"

#flag -lcsfml-graphics
