module window

// WindowHandle: low-level window handle type
pub type WindowHandle = voidptr
