// network: socket-based communication, utilities and higher-level network protocols (HTTP, FTP)
module network

#flag -lcsfml-network