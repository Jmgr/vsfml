module network

#include <SFML/Network/Export.h>
