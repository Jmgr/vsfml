module system

#include <SFML/System/Export.h>
