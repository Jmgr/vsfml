module graphics

// color_black: black predefined color
pub const color_black = color_from_rgb(0, 0, 0)

// color_white: white predefined color
pub const color_white = color_from_rgb(255, 255, 255)

// color_red: red predefined color
pub const color_red = color_from_rgb(255, 0, 0)

// color_green: green predefined color
pub const color_green = color_from_rgb(0, 255, 0)

// color_blue: blue predefined color
pub const color_blue = color_from_rgb(0, 0, 255)

// color_yellow: yellow predefined color
pub const color_yellow = color_from_rgb(255, 255, 0)

// color_magenta: magenta predefined color
pub const color_magenta = color_from_rgb(255, 0, 255)

// color_cyan: cyan predefined color
pub const color_cyan = color_from_rgb(0, 255, 255)

// color_transparent: transparent (black) predefined color
pub const color_transparent = color_from_rgba(0, 0, 0, 0)
