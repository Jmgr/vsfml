module graphics

#include <SFML/Graphics/Export.h>
