module graphics

#include <SFML/Graphics/Types.h>

struct C.sfCircleShape {
}

// CircleShape
pub type CircleShape = C.sfCircleShape

struct C.sfConvexShape {
}

// ConvexShape
pub type ConvexShape = C.sfConvexShape

struct C.sfFont {
}

// Font
pub type Font = C.sfFont

struct C.sfImage {
}

// Image
pub type Image = C.sfImage

struct C.sfShader {
}

// Shader
pub type Shader = C.sfShader

struct C.sfRectangleShape {
}

// RectangleShape
pub type RectangleShape = C.sfRectangleShape

struct C.sfRenderTexture {
}

// RenderTexture
pub type RenderTexture = C.sfRenderTexture

struct C.sfRenderWindow {
}

// RenderWindow
pub type RenderWindow = C.sfRenderWindow

struct C.sfShape {
}

// Shape
pub type Shape = C.sfShape

struct C.sfSprite {
}

// Sprite
pub type Sprite = C.sfSprite

struct C.sfText {
}

// Text
pub type Text = C.sfText

struct C.sfTexture {
}

// Texture
pub type Texture = C.sfTexture

struct C.sfTransformable {
}

// Transformable
pub type Transformable = C.sfTransformable

struct C.sfVertexArray {
}

// VertexArray
pub type VertexArray = C.sfVertexArray

struct C.sfVertexBuffer {
}

// VertexBuffer
pub type VertexBuffer = C.sfVertexBuffer

struct C.sfView {
}

// View
pub type View = C.sfView
