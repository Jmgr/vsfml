// Copyright(C) 2021 Jonathan Mercier-Ganady
// For conditions of distribution and use, see the LICENSE file

module vsfml
