module audio

#include <SFML/Audio/Export.h>
